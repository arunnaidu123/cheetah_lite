LIBRARY ieee;
USE ieee.std_logic_1164.all;

TYPE fortyeight IS RECORD
	test : STD_LOGIC_VECTOR(48-1 DOWNTO 0);
END RECORD;

